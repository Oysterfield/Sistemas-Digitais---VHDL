library ieee;
use ieee.std_logic_1164.all;


entity AcessoARAM is
	port(
	);
end entity;

architecture estrutura os AcessoARAM is
begin
end;